localparam  RV32_OPC_DET = 2'b11;
localparam  RV32_OPC_B = 5'b11000;
localparam  RV32_OPC_JALR = 5'b11001;
localparam  RV32_OPC_JAL = 5'b11011;
