`define SLAVE_SEL_WIDTH                 4
`define TCM_ADDR_WIDTH                  11

`define BRANCH_PREDICTION_SIMPLE
