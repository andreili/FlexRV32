typedef struct packed
{
} wb_bus_t;
